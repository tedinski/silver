grammar silver_features:anno_short_names:c;

synthesized attribute foo :: String;
