grammar silver_features:anno_short_names:b;

annotation foo :: String;
synthesized attribute baz :: String;
