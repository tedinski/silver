grammar silver_features:anno_short_names:a;

annotation foo :: String;
synthesized attribute baz :: String;