grammar silver:compiler:extension:opersection;

imports silver:compiler:definition:core;
imports silver:compiler:definition:type:syntax;
imports silver:compiler:definition:type;

imports silver:compiler:metatranslation;

imports silver:compiler:extension:silverconstruction;